-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb0",
     9 => x"8c080b0b",
    10 => x"0bb09008",
    11 => x"0b0b0bb0",
    12 => x"94080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b0940c0b",
    16 => x"0b0bb090",
    17 => x"0c0b0b0b",
    18 => x"b08c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba880",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b08c70b5",
    57 => x"b0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"88c40402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"b09c0c9f",
    65 => x"0bb0a00c",
    66 => x"a0717081",
    67 => x"055334b0",
    68 => x"a008ff05",
    69 => x"b0a00cb0",
    70 => x"a0088025",
    71 => x"eb38b09c",
    72 => x"08ff05b0",
    73 => x"9c0cb09c",
    74 => x"088025d7",
    75 => x"38800bb0",
    76 => x"a00c800b",
    77 => x"b09c0c02",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"b09c0825",
    97 => x"8f3882bc",
    98 => x"2db09c08",
    99 => x"ff05b09c",
   100 => x"0c82fe04",
   101 => x"b09c08b0",
   102 => x"a0085351",
   103 => x"728a2e09",
   104 => x"8106b738",
   105 => x"7151719f",
   106 => x"24a038b0",
   107 => x"9c08a029",
   108 => x"11f88011",
   109 => x"5151a071",
   110 => x"34b0a008",
   111 => x"8105b0a0",
   112 => x"0cb0a008",
   113 => x"519f7125",
   114 => x"e238800b",
   115 => x"b0a00cb0",
   116 => x"9c088105",
   117 => x"b09c0c83",
   118 => x"ee0470a0",
   119 => x"2912f880",
   120 => x"11515172",
   121 => x"7134b0a0",
   122 => x"088105b0",
   123 => x"a00cb0a0",
   124 => x"08a02e09",
   125 => x"81068e38",
   126 => x"800bb0a0",
   127 => x"0cb09c08",
   128 => x"8105b09c",
   129 => x"0c028c05",
   130 => x"0d0402e8",
   131 => x"050d7779",
   132 => x"5656880b",
   133 => x"fc167771",
   134 => x"2c8f0654",
   135 => x"52548053",
   136 => x"72722595",
   137 => x"387153fb",
   138 => x"e0145187",
   139 => x"71348114",
   140 => x"ff145454",
   141 => x"72f13871",
   142 => x"53f91576",
   143 => x"712c8706",
   144 => x"53517180",
   145 => x"2e8b38fb",
   146 => x"e0145171",
   147 => x"71348114",
   148 => x"54728e24",
   149 => x"95388f73",
   150 => x"3153fbe0",
   151 => x"1451a071",
   152 => x"348114ff",
   153 => x"14545472",
   154 => x"f1380298",
   155 => x"050d0402",
   156 => x"ec050d80",
   157 => x"0bb0a40c",
   158 => x"f68c08f6",
   159 => x"90087188",
   160 => x"2c565481",
   161 => x"ff065273",
   162 => x"72258838",
   163 => x"7154820b",
   164 => x"b0a40c72",
   165 => x"882c7381",
   166 => x"ff065455",
   167 => x"7473258b",
   168 => x"3872b0a4",
   169 => x"088407b0",
   170 => x"a40c5573",
   171 => x"842b86a0",
   172 => x"71258371",
   173 => x"31700b0b",
   174 => x"0bad900c",
   175 => x"81712bff",
   176 => x"05f6880c",
   177 => x"fdfc13ff",
   178 => x"122c7888",
   179 => x"29ff9405",
   180 => x"70812cb0",
   181 => x"a4085258",
   182 => x"52555152",
   183 => x"5476802e",
   184 => x"85387081",
   185 => x"075170f6",
   186 => x"940c7109",
   187 => x"8105f680",
   188 => x"0c720981",
   189 => x"05f6840c",
   190 => x"0294050d",
   191 => x"0402f405",
   192 => x"0d745372",
   193 => x"70810554",
   194 => x"80f52d52",
   195 => x"71802e89",
   196 => x"38715182",
   197 => x"f82d8683",
   198 => x"04810bb0",
   199 => x"8c0c028c",
   200 => x"050d0402",
   201 => x"fc050d81",
   202 => x"808051c0",
   203 => x"115170fb",
   204 => x"38028405",
   205 => x"0d0402fc",
   206 => x"050d84bf",
   207 => x"5186a32d",
   208 => x"ff115170",
   209 => x"8025f638",
   210 => x"0284050d",
   211 => x"0402fc05",
   212 => x"0dec5183",
   213 => x"710c86a3",
   214 => x"2d82710c",
   215 => x"0284050d",
   216 => x"0402fc05",
   217 => x"0dec5192",
   218 => x"710c86a3",
   219 => x"2d82710c",
   220 => x"0284050d",
   221 => x"0402dc05",
   222 => x"0d7a5480",
   223 => x"7453b0a8",
   224 => x"5259a4d2",
   225 => x"2db08c08",
   226 => x"792e8191",
   227 => x"38b0ac08",
   228 => x"70f80c89",
   229 => x"1580f52d",
   230 => x"8a1680f5",
   231 => x"2d718280",
   232 => x"29058817",
   233 => x"80f52d70",
   234 => x"84808029",
   235 => x"12f40c57",
   236 => x"555755a4",
   237 => x"0bec0c78",
   238 => x"ff165558",
   239 => x"73792e8b",
   240 => x"38811874",
   241 => x"812a5558",
   242 => x"73f738f7",
   243 => x"18588159",
   244 => x"80752580",
   245 => x"c8387752",
   246 => x"7351848a",
   247 => x"2db0f452",
   248 => x"b0a851a7",
   249 => x"882db08c",
   250 => x"08802e9a",
   251 => x"38b0f457",
   252 => x"83fc5676",
   253 => x"70840558",
   254 => x"08e80cfc",
   255 => x"16567580",
   256 => x"25f13888",
   257 => x"8d04b08c",
   258 => x"08598480",
   259 => x"55b0a851",
   260 => x"a6db2dfc",
   261 => x"80158115",
   262 => x"555587d0",
   263 => x"0486b62d",
   264 => x"840bec0c",
   265 => x"78802e8d",
   266 => x"38ad9451",
   267 => x"8fe22d8d",
   268 => x"e52d88bb",
   269 => x"04af9851",
   270 => x"8fe22d78",
   271 => x"b08c0c02",
   272 => x"a4050d04",
   273 => x"02ec050d",
   274 => x"840bec0c",
   275 => x"8dcd2d8a",
   276 => x"b72d81f7",
   277 => x"2d9ea12d",
   278 => x"b08c0880",
   279 => x"2e81c338",
   280 => x"86f551a7",
   281 => x"fa2dad94",
   282 => x"518fe22d",
   283 => x"8de52d8a",
   284 => x"c32d8ff2",
   285 => x"2dadc00b",
   286 => x"80f52d70",
   287 => x"8a2b9880",
   288 => x"06adcc0b",
   289 => x"80f52d70",
   290 => x"8c2ba080",
   291 => x"06add80b",
   292 => x"80f52d70",
   293 => x"822b8406",
   294 => x"74730707",
   295 => x"ade40b80",
   296 => x"f52d708d",
   297 => x"2b80c080",
   298 => x"06adf00b",
   299 => x"80f52d70",
   300 => x"832b8806",
   301 => x"74730707",
   302 => x"adfc0b80",
   303 => x"f52d7084",
   304 => x"2bb006ae",
   305 => x"880b80f5",
   306 => x"2d70862b",
   307 => x"80c00674",
   308 => x"730707ae",
   309 => x"940b80f5",
   310 => x"2d70872b",
   311 => x"818006ae",
   312 => x"a00b80f5",
   313 => x"2d70892b",
   314 => x"84800674",
   315 => x"730707ae",
   316 => x"ac0b80f5",
   317 => x"2d708e2b",
   318 => x"83808006",
   319 => x"7207fc0c",
   320 => x"53545454",
   321 => x"54545454",
   322 => x"54545454",
   323 => x"56545257",
   324 => x"57535386",
   325 => x"52b08c08",
   326 => x"83388452",
   327 => x"71ec0c88",
   328 => x"ef04800b",
   329 => x"b08c0c02",
   330 => x"94050d04",
   331 => x"71980c04",
   332 => x"ffb008b0",
   333 => x"8c0c0481",
   334 => x"0bffb00c",
   335 => x"04800bff",
   336 => x"b00c0402",
   337 => x"f4050d8b",
   338 => x"c504b08c",
   339 => x"0881f02e",
   340 => x"09810689",
   341 => x"38810baf",
   342 => x"fc0c8bc5",
   343 => x"04b08c08",
   344 => x"81e02e09",
   345 => x"81068938",
   346 => x"810bb080",
   347 => x"0c8bc504",
   348 => x"b08c0852",
   349 => x"b0800880",
   350 => x"2e8838b0",
   351 => x"8c088180",
   352 => x"05527184",
   353 => x"2c728f06",
   354 => x"5353affc",
   355 => x"08802e99",
   356 => x"38728429",
   357 => x"afbc0572",
   358 => x"1381712b",
   359 => x"70097308",
   360 => x"06730c51",
   361 => x"53538bbb",
   362 => x"04728429",
   363 => x"afbc0572",
   364 => x"1383712b",
   365 => x"72080772",
   366 => x"0c535380",
   367 => x"0bb0800c",
   368 => x"800baffc",
   369 => x"0cb0b451",
   370 => x"8cc62db0",
   371 => x"8c08ff24",
   372 => x"fef83880",
   373 => x"0bb08c0c",
   374 => x"028c050d",
   375 => x"0402f805",
   376 => x"0dafbc52",
   377 => x"8f518072",
   378 => x"70840554",
   379 => x"0cff1151",
   380 => x"708025f2",
   381 => x"38028805",
   382 => x"0d0402f0",
   383 => x"050d7551",
   384 => x"8abd2d70",
   385 => x"822cfc06",
   386 => x"afbc1172",
   387 => x"109e0671",
   388 => x"0870722a",
   389 => x"70830682",
   390 => x"742b7009",
   391 => x"7406760c",
   392 => x"54515657",
   393 => x"5351538a",
   394 => x"b72d71b0",
   395 => x"8c0c0290",
   396 => x"050d0402",
   397 => x"fc050d72",
   398 => x"5180710c",
   399 => x"800b8412",
   400 => x"0c028405",
   401 => x"0d0402f0",
   402 => x"050d7570",
   403 => x"08841208",
   404 => x"535353ff",
   405 => x"5471712e",
   406 => x"a8388abd",
   407 => x"2d841308",
   408 => x"70842914",
   409 => x"88117008",
   410 => x"7081ff06",
   411 => x"84180881",
   412 => x"11870684",
   413 => x"1a0c5351",
   414 => x"55515151",
   415 => x"8ab72d71",
   416 => x"5473b08c",
   417 => x"0c029005",
   418 => x"0d0402f8",
   419 => x"050d8abd",
   420 => x"2de00870",
   421 => x"8b2a7081",
   422 => x"06515252",
   423 => x"70802e9d",
   424 => x"38b0b408",
   425 => x"708429b0",
   426 => x"bc057381",
   427 => x"ff06710c",
   428 => x"5151b0b4",
   429 => x"08811187",
   430 => x"06b0b40c",
   431 => x"51800bb0",
   432 => x"dc0c8ab0",
   433 => x"2d8ab72d",
   434 => x"0288050d",
   435 => x"0402fc05",
   436 => x"0db0b451",
   437 => x"8cb32d8b",
   438 => x"dd2d8d8a",
   439 => x"518aac2d",
   440 => x"0284050d",
   441 => x"0402fc05",
   442 => x"0d8def04",
   443 => x"8ac32d80",
   444 => x"f6518bfa",
   445 => x"2db08c08",
   446 => x"f33880da",
   447 => x"518bfa2d",
   448 => x"b08c08e8",
   449 => x"38b08c08",
   450 => x"b0880cb0",
   451 => x"8c085184",
   452 => x"ef2d0284",
   453 => x"050d0402",
   454 => x"ec050d76",
   455 => x"54805287",
   456 => x"0b881580",
   457 => x"f52d5653",
   458 => x"74722483",
   459 => x"38a05372",
   460 => x"5182f82d",
   461 => x"81128b15",
   462 => x"80f52d54",
   463 => x"52727225",
   464 => x"de380294",
   465 => x"050d0402",
   466 => x"f0050db0",
   467 => x"e0085481",
   468 => x"f72d800b",
   469 => x"b0e40c73",
   470 => x"08802e81",
   471 => x"8038820b",
   472 => x"b0a00cb0",
   473 => x"e4088f06",
   474 => x"b09c0c73",
   475 => x"08527183",
   476 => x"2e963871",
   477 => x"83268938",
   478 => x"71812eaf",
   479 => x"388fc804",
   480 => x"71852e9f",
   481 => x"388fc804",
   482 => x"881480f5",
   483 => x"2d841508",
   484 => x"abe45354",
   485 => x"5285fd2d",
   486 => x"71842913",
   487 => x"70085252",
   488 => x"8fcc0473",
   489 => x"518e972d",
   490 => x"8fc804b0",
   491 => x"84088815",
   492 => x"082c7081",
   493 => x"06515271",
   494 => x"802e8738",
   495 => x"abe8518f",
   496 => x"c504abec",
   497 => x"5185fd2d",
   498 => x"84140851",
   499 => x"85fd2db0",
   500 => x"e4088105",
   501 => x"b0e40c8c",
   502 => x"14548ed7",
   503 => x"04029005",
   504 => x"0d0471b0",
   505 => x"e00c8ec7",
   506 => x"2db0e408",
   507 => x"ff05b0e8",
   508 => x"0c0402e8",
   509 => x"050db0e0",
   510 => x"08b0ec08",
   511 => x"57558751",
   512 => x"8bfa2db0",
   513 => x"8c08812a",
   514 => x"70810651",
   515 => x"5271802e",
   516 => x"a0389098",
   517 => x"048ac32d",
   518 => x"87518bfa",
   519 => x"2db08c08",
   520 => x"f438b088",
   521 => x"08813270",
   522 => x"b0880c70",
   523 => x"525284ef",
   524 => x"2d80fe51",
   525 => x"8bfa2db0",
   526 => x"8c08802e",
   527 => x"a638b088",
   528 => x"08802e91",
   529 => x"38800bb0",
   530 => x"880c8051",
   531 => x"84ef2d90",
   532 => x"d5048ac3",
   533 => x"2d80fe51",
   534 => x"8bfa2db0",
   535 => x"8c08f338",
   536 => x"86e12db0",
   537 => x"88089038",
   538 => x"81fd518b",
   539 => x"fa2d81fa",
   540 => x"518bfa2d",
   541 => x"96a80481",
   542 => x"f5518bfa",
   543 => x"2db08c08",
   544 => x"812a7081",
   545 => x"06515271",
   546 => x"802eaf38",
   547 => x"b0e80852",
   548 => x"71802e89",
   549 => x"38ff12b0",
   550 => x"e80c91ba",
   551 => x"04b0e408",
   552 => x"10b0e408",
   553 => x"05708429",
   554 => x"16515288",
   555 => x"1208802e",
   556 => x"8938ff51",
   557 => x"88120852",
   558 => x"712d81f2",
   559 => x"518bfa2d",
   560 => x"b08c0881",
   561 => x"2a708106",
   562 => x"51527180",
   563 => x"2eb138b0",
   564 => x"e408ff11",
   565 => x"b0e80856",
   566 => x"53537372",
   567 => x"25893881",
   568 => x"14b0e80c",
   569 => x"91ff0472",
   570 => x"10137084",
   571 => x"29165152",
   572 => x"88120880",
   573 => x"2e8938fe",
   574 => x"51881208",
   575 => x"52712d81",
   576 => x"fd518bfa",
   577 => x"2db08c08",
   578 => x"812a7081",
   579 => x"06515271",
   580 => x"802ead38",
   581 => x"b0e80880",
   582 => x"2e893880",
   583 => x"0bb0e80c",
   584 => x"92c004b0",
   585 => x"e40810b0",
   586 => x"e4080570",
   587 => x"84291651",
   588 => x"52881208",
   589 => x"802e8938",
   590 => x"fd518812",
   591 => x"0852712d",
   592 => x"81fa518b",
   593 => x"fa2db08c",
   594 => x"08812a70",
   595 => x"81065152",
   596 => x"71802eae",
   597 => x"38b0e408",
   598 => x"ff115452",
   599 => x"b0e80873",
   600 => x"25883872",
   601 => x"b0e80c93",
   602 => x"82047110",
   603 => x"12708429",
   604 => x"16515288",
   605 => x"1208802e",
   606 => x"8938fc51",
   607 => x"88120852",
   608 => x"712db0e8",
   609 => x"08705354",
   610 => x"73802e8a",
   611 => x"388c15ff",
   612 => x"15555593",
   613 => x"8804820b",
   614 => x"b0a00c71",
   615 => x"8f06b09c",
   616 => x"0c81eb51",
   617 => x"8bfa2db0",
   618 => x"8c08812a",
   619 => x"70810651",
   620 => x"5271802e",
   621 => x"ad387408",
   622 => x"852e0981",
   623 => x"06a43888",
   624 => x"1580f52d",
   625 => x"ff055271",
   626 => x"881681b7",
   627 => x"2d71982b",
   628 => x"52718025",
   629 => x"8838800b",
   630 => x"881681b7",
   631 => x"2d74518e",
   632 => x"972d81f4",
   633 => x"518bfa2d",
   634 => x"b08c0881",
   635 => x"2a708106",
   636 => x"51527180",
   637 => x"2eb33874",
   638 => x"08852e09",
   639 => x"8106aa38",
   640 => x"881580f5",
   641 => x"2d810552",
   642 => x"71881681",
   643 => x"b72d7181",
   644 => x"ff068b16",
   645 => x"80f52d54",
   646 => x"52727227",
   647 => x"87387288",
   648 => x"1681b72d",
   649 => x"74518e97",
   650 => x"2d80da51",
   651 => x"8bfa2db0",
   652 => x"8c08812a",
   653 => x"70810651",
   654 => x"5271802e",
   655 => x"81a638b0",
   656 => x"e008b0e8",
   657 => x"08555373",
   658 => x"802e8a38",
   659 => x"8c13ff15",
   660 => x"555394c7",
   661 => x"04720852",
   662 => x"71822ea6",
   663 => x"38718226",
   664 => x"89387181",
   665 => x"2ea93895",
   666 => x"e4047183",
   667 => x"2eb13871",
   668 => x"842e0981",
   669 => x"0680ed38",
   670 => x"88130851",
   671 => x"8fe22d95",
   672 => x"e404b0e8",
   673 => x"08518813",
   674 => x"0852712d",
   675 => x"95e40481",
   676 => x"0b881408",
   677 => x"2bb08408",
   678 => x"32b0840c",
   679 => x"95ba0488",
   680 => x"1380f52d",
   681 => x"81058b14",
   682 => x"80f52d53",
   683 => x"54717424",
   684 => x"83388054",
   685 => x"73881481",
   686 => x"b72d8ec7",
   687 => x"2d95e404",
   688 => x"7508802e",
   689 => x"a2387508",
   690 => x"518bfa2d",
   691 => x"b08c0881",
   692 => x"06527180",
   693 => x"2e8b38b0",
   694 => x"e8085184",
   695 => x"16085271",
   696 => x"2d881656",
   697 => x"75da3880",
   698 => x"54800bb0",
   699 => x"a00c738f",
   700 => x"06b09c0c",
   701 => x"a05273b0",
   702 => x"e8082e09",
   703 => x"81069838",
   704 => x"b0e408ff",
   705 => x"05743270",
   706 => x"09810570",
   707 => x"72079f2a",
   708 => x"91713151",
   709 => x"51535371",
   710 => x"5182f82d",
   711 => x"8114548e",
   712 => x"7425c638",
   713 => x"b0880852",
   714 => x"71b08c0c",
   715 => x"0298050d",
   716 => x"0402f405",
   717 => x"0dd45281",
   718 => x"ff720c71",
   719 => x"085381ff",
   720 => x"720c7288",
   721 => x"2b83fe80",
   722 => x"06720870",
   723 => x"81ff0651",
   724 => x"525381ff",
   725 => x"720c7271",
   726 => x"07882b72",
   727 => x"087081ff",
   728 => x"06515253",
   729 => x"81ff720c",
   730 => x"72710788",
   731 => x"2b720870",
   732 => x"81ff0672",
   733 => x"07b08c0c",
   734 => x"5253028c",
   735 => x"050d0402",
   736 => x"f4050d74",
   737 => x"767181ff",
   738 => x"06d40c53",
   739 => x"53b0f008",
   740 => x"85387189",
   741 => x"2b527198",
   742 => x"2ad40c71",
   743 => x"902a7081",
   744 => x"ff06d40c",
   745 => x"5171882a",
   746 => x"7081ff06",
   747 => x"d40c5171",
   748 => x"81ff06d4",
   749 => x"0c72902a",
   750 => x"7081ff06",
   751 => x"d40c51d4",
   752 => x"087081ff",
   753 => x"06515182",
   754 => x"b8bf5270",
   755 => x"81ff2e09",
   756 => x"81069438",
   757 => x"81ff0bd4",
   758 => x"0cd40870",
   759 => x"81ff06ff",
   760 => x"14545151",
   761 => x"71e53870",
   762 => x"b08c0c02",
   763 => x"8c050d04",
   764 => x"02fc050d",
   765 => x"81c75181",
   766 => x"ff0bd40c",
   767 => x"ff115170",
   768 => x"8025f438",
   769 => x"0284050d",
   770 => x"0402f405",
   771 => x"0d81ff0b",
   772 => x"d40c9353",
   773 => x"805287fc",
   774 => x"80c15196",
   775 => x"ff2db08c",
   776 => x"088b3881",
   777 => x"ff0bd40c",
   778 => x"815398b6",
   779 => x"0497f02d",
   780 => x"ff135372",
   781 => x"df3872b0",
   782 => x"8c0c028c",
   783 => x"050d0402",
   784 => x"ec050d81",
   785 => x"0bb0f00c",
   786 => x"8454d008",
   787 => x"708f2a70",
   788 => x"81065151",
   789 => x"5372f338",
   790 => x"72d00c97",
   791 => x"f02dabf0",
   792 => x"5185fd2d",
   793 => x"d008708f",
   794 => x"2a708106",
   795 => x"51515372",
   796 => x"f338810b",
   797 => x"d00cb153",
   798 => x"805284d4",
   799 => x"80c05196",
   800 => x"ff2db08c",
   801 => x"08812e93",
   802 => x"3872822e",
   803 => x"bd38ff13",
   804 => x"5372e538",
   805 => x"ff145473",
   806 => x"ffb03897",
   807 => x"f02d83aa",
   808 => x"52849c80",
   809 => x"c85196ff",
   810 => x"2db08c08",
   811 => x"812e0981",
   812 => x"06923896",
   813 => x"b12db08c",
   814 => x"0883ffff",
   815 => x"06537283",
   816 => x"aa2e9d38",
   817 => x"98892d99",
   818 => x"db04abfc",
   819 => x"5185fd2d",
   820 => x"80539ba9",
   821 => x"04ac9451",
   822 => x"85fd2d80",
   823 => x"549afb04",
   824 => x"81ff0bd4",
   825 => x"0cb15497",
   826 => x"f02d8fcf",
   827 => x"53805287",
   828 => x"fc80f751",
   829 => x"96ff2db0",
   830 => x"8c0855b0",
   831 => x"8c08812e",
   832 => x"0981069b",
   833 => x"3881ff0b",
   834 => x"d40c820a",
   835 => x"52849c80",
   836 => x"e95196ff",
   837 => x"2db08c08",
   838 => x"802e8d38",
   839 => x"97f02dff",
   840 => x"135372c9",
   841 => x"389aee04",
   842 => x"81ff0bd4",
   843 => x"0cb08c08",
   844 => x"5287fc80",
   845 => x"fa5196ff",
   846 => x"2db08c08",
   847 => x"b13881ff",
   848 => x"0bd40cd4",
   849 => x"085381ff",
   850 => x"0bd40c81",
   851 => x"ff0bd40c",
   852 => x"81ff0bd4",
   853 => x"0c81ff0b",
   854 => x"d40c7286",
   855 => x"2a708106",
   856 => x"76565153",
   857 => x"729538b0",
   858 => x"8c08549a",
   859 => x"fb047382",
   860 => x"2efee238",
   861 => x"ff145473",
   862 => x"feed3873",
   863 => x"b0f00c73",
   864 => x"8b388152",
   865 => x"87fc80d0",
   866 => x"5196ff2d",
   867 => x"81ff0bd4",
   868 => x"0cd00870",
   869 => x"8f2a7081",
   870 => x"06515153",
   871 => x"72f33872",
   872 => x"d00c81ff",
   873 => x"0bd40c81",
   874 => x"5372b08c",
   875 => x"0c029405",
   876 => x"0d0402e8",
   877 => x"050d7855",
   878 => x"805681ff",
   879 => x"0bd40cd0",
   880 => x"08708f2a",
   881 => x"70810651",
   882 => x"515372f3",
   883 => x"3882810b",
   884 => x"d00c81ff",
   885 => x"0bd40c77",
   886 => x"5287fc80",
   887 => x"d15196ff",
   888 => x"2d80dbc6",
   889 => x"df54b08c",
   890 => x"08802e8a",
   891 => x"38acb451",
   892 => x"85fd2d9c",
   893 => x"c90481ff",
   894 => x"0bd40cd4",
   895 => x"087081ff",
   896 => x"06515372",
   897 => x"81fe2e09",
   898 => x"81069d38",
   899 => x"80ff5396",
   900 => x"b12db08c",
   901 => x"08757084",
   902 => x"05570cff",
   903 => x"13537280",
   904 => x"25ed3881",
   905 => x"569cae04",
   906 => x"ff145473",
   907 => x"c93881ff",
   908 => x"0bd40c81",
   909 => x"ff0bd40c",
   910 => x"d008708f",
   911 => x"2a708106",
   912 => x"51515372",
   913 => x"f33872d0",
   914 => x"0c75b08c",
   915 => x"0c029805",
   916 => x"0d0402e8",
   917 => x"050d7779",
   918 => x"7b585555",
   919 => x"80537276",
   920 => x"25a33874",
   921 => x"70810556",
   922 => x"80f52d74",
   923 => x"70810556",
   924 => x"80f52d52",
   925 => x"5271712e",
   926 => x"86388151",
   927 => x"9d870481",
   928 => x"13539cde",
   929 => x"04805170",
   930 => x"b08c0c02",
   931 => x"98050d04",
   932 => x"02ec050d",
   933 => x"76557480",
   934 => x"2ebb389a",
   935 => x"1580e02d",
   936 => x"51a7de2d",
   937 => x"b08c08b0",
   938 => x"8c08b5a0",
   939 => x"0cb08c08",
   940 => x"5454b4fc",
   941 => x"08802e99",
   942 => x"38941580",
   943 => x"e02d51a7",
   944 => x"de2db08c",
   945 => x"08902b83",
   946 => x"fff00a06",
   947 => x"70750751",
   948 => x"5372b5a0",
   949 => x"0cb5a008",
   950 => x"5372802e",
   951 => x"9938b4f4",
   952 => x"08fe1471",
   953 => x"29b58808",
   954 => x"05b5a40c",
   955 => x"70842bb5",
   956 => x"800c549e",
   957 => x"9c04b58c",
   958 => x"08b5a00c",
   959 => x"b59008b5",
   960 => x"a40cb4fc",
   961 => x"08802e8a",
   962 => x"38b4f408",
   963 => x"842b539e",
   964 => x"9804b594",
   965 => x"08842b53",
   966 => x"72b5800c",
   967 => x"0294050d",
   968 => x"0402d805",
   969 => x"0d800bb4",
   970 => x"fc0c8454",
   971 => x"98bf2db0",
   972 => x"8c08802e",
   973 => x"9538b0f4",
   974 => x"5280519b",
   975 => x"b22db08c",
   976 => x"08802e86",
   977 => x"38fe549e",
   978 => x"d204ff14",
   979 => x"54738024",
   980 => x"db38738c",
   981 => x"38acc451",
   982 => x"85fd2d73",
   983 => x"55a3db04",
   984 => x"8056810b",
   985 => x"b5a80c88",
   986 => x"53acd852",
   987 => x"b1aa519c",
   988 => x"d22db08c",
   989 => x"08762e09",
   990 => x"81068738",
   991 => x"b08c08b5",
   992 => x"a80c8853",
   993 => x"ace452b1",
   994 => x"c6519cd2",
   995 => x"2db08c08",
   996 => x"8738b08c",
   997 => x"08b5a80c",
   998 => x"b5a80880",
   999 => x"2e80f638",
  1000 => x"b4ba0b80",
  1001 => x"f52db4bb",
  1002 => x"0b80f52d",
  1003 => x"71982b71",
  1004 => x"902b07b4",
  1005 => x"bc0b80f5",
  1006 => x"2d70882b",
  1007 => x"7207b4bd",
  1008 => x"0b80f52d",
  1009 => x"7107b4f2",
  1010 => x"0b80f52d",
  1011 => x"b4f30b80",
  1012 => x"f52d7188",
  1013 => x"2b07535f",
  1014 => x"54525a56",
  1015 => x"57557381",
  1016 => x"abaa2e09",
  1017 => x"81068d38",
  1018 => x"7551a7ae",
  1019 => x"2db08c08",
  1020 => x"56a08104",
  1021 => x"7382d4d5",
  1022 => x"2e8738ac",
  1023 => x"f051a0c2",
  1024 => x"04b0f452",
  1025 => x"75519bb2",
  1026 => x"2db08c08",
  1027 => x"55b08c08",
  1028 => x"802e83c7",
  1029 => x"388853ac",
  1030 => x"e452b1c6",
  1031 => x"519cd22d",
  1032 => x"b08c0889",
  1033 => x"38810bb4",
  1034 => x"fc0ca0c8",
  1035 => x"048853ac",
  1036 => x"d852b1aa",
  1037 => x"519cd22d",
  1038 => x"b08c0880",
  1039 => x"2e8a38ad",
  1040 => x"845185fd",
  1041 => x"2da1a204",
  1042 => x"b4f20b80",
  1043 => x"f52d5473",
  1044 => x"80d52e09",
  1045 => x"810680ca",
  1046 => x"38b4f30b",
  1047 => x"80f52d54",
  1048 => x"7381aa2e",
  1049 => x"098106ba",
  1050 => x"38800bb0",
  1051 => x"f40b80f5",
  1052 => x"2d565474",
  1053 => x"81e92e83",
  1054 => x"38815474",
  1055 => x"81eb2e8c",
  1056 => x"38805573",
  1057 => x"752e0981",
  1058 => x"0682d038",
  1059 => x"b0ff0b80",
  1060 => x"f52d5574",
  1061 => x"8d38b180",
  1062 => x"0b80f52d",
  1063 => x"5473822e",
  1064 => x"86388055",
  1065 => x"a3db04b1",
  1066 => x"810b80f5",
  1067 => x"2d70b4f4",
  1068 => x"0cff05b4",
  1069 => x"f80cb182",
  1070 => x"0b80f52d",
  1071 => x"b1830b80",
  1072 => x"f52d5876",
  1073 => x"05778280",
  1074 => x"290570b5",
  1075 => x"840cb184",
  1076 => x"0b80f52d",
  1077 => x"70b5980c",
  1078 => x"b4fc0859",
  1079 => x"57587680",
  1080 => x"2e81a338",
  1081 => x"8853ace4",
  1082 => x"52b1c651",
  1083 => x"9cd22db0",
  1084 => x"8c0881e7",
  1085 => x"38b4f408",
  1086 => x"70842bb5",
  1087 => x"800c70b5",
  1088 => x"940cb199",
  1089 => x"0b80f52d",
  1090 => x"b1980b80",
  1091 => x"f52d7182",
  1092 => x"802905b1",
  1093 => x"9a0b80f5",
  1094 => x"2d708480",
  1095 => x"802912b1",
  1096 => x"9b0b80f5",
  1097 => x"2d708180",
  1098 => x"0a291270",
  1099 => x"b59c0cb5",
  1100 => x"98087129",
  1101 => x"b5840805",
  1102 => x"70b5880c",
  1103 => x"b1a10b80",
  1104 => x"f52db1a0",
  1105 => x"0b80f52d",
  1106 => x"71828029",
  1107 => x"05b1a20b",
  1108 => x"80f52d70",
  1109 => x"84808029",
  1110 => x"12b1a30b",
  1111 => x"80f52d70",
  1112 => x"982b81f0",
  1113 => x"0a067205",
  1114 => x"70b58c0c",
  1115 => x"fe117e29",
  1116 => x"7705b590",
  1117 => x"0c525952",
  1118 => x"43545e51",
  1119 => x"5259525d",
  1120 => x"575957a3",
  1121 => x"d404b186",
  1122 => x"0b80f52d",
  1123 => x"b1850b80",
  1124 => x"f52d7182",
  1125 => x"80290570",
  1126 => x"b5800c70",
  1127 => x"a02983ff",
  1128 => x"0570892a",
  1129 => x"70b5940c",
  1130 => x"b18b0b80",
  1131 => x"f52db18a",
  1132 => x"0b80f52d",
  1133 => x"71828029",
  1134 => x"0570b59c",
  1135 => x"0c7b7129",
  1136 => x"1e70b590",
  1137 => x"0c7db58c",
  1138 => x"0c7305b5",
  1139 => x"880c555e",
  1140 => x"51515555",
  1141 => x"80519d90",
  1142 => x"2d815574",
  1143 => x"b08c0c02",
  1144 => x"a8050d04",
  1145 => x"02ec050d",
  1146 => x"7670872c",
  1147 => x"7180ff06",
  1148 => x"555654b4",
  1149 => x"fc088a38",
  1150 => x"73882c74",
  1151 => x"81ff0654",
  1152 => x"55b0f452",
  1153 => x"b5840815",
  1154 => x"519bb22d",
  1155 => x"b08c0854",
  1156 => x"b08c0880",
  1157 => x"2eb338b4",
  1158 => x"fc08802e",
  1159 => x"98387284",
  1160 => x"29b0f405",
  1161 => x"70085253",
  1162 => x"a7ae2db0",
  1163 => x"8c08f00a",
  1164 => x"0653a4c7",
  1165 => x"047210b0",
  1166 => x"f4057080",
  1167 => x"e02d5253",
  1168 => x"a7de2db0",
  1169 => x"8c085372",
  1170 => x"5473b08c",
  1171 => x"0c029405",
  1172 => x"0d0402cc",
  1173 => x"050d7e60",
  1174 => x"5e5a800b",
  1175 => x"b5a008b5",
  1176 => x"a408595c",
  1177 => x"568058b5",
  1178 => x"8008782e",
  1179 => x"81ae3877",
  1180 => x"8f06a017",
  1181 => x"5754738f",
  1182 => x"38b0f452",
  1183 => x"76518117",
  1184 => x"579bb22d",
  1185 => x"b0f45680",
  1186 => x"7680f52d",
  1187 => x"56547474",
  1188 => x"2e833881",
  1189 => x"547481e5",
  1190 => x"2e80f638",
  1191 => x"81707506",
  1192 => x"555c7380",
  1193 => x"2e80ea38",
  1194 => x"8b1680f5",
  1195 => x"2d980659",
  1196 => x"7880de38",
  1197 => x"8b537c52",
  1198 => x"75519cd2",
  1199 => x"2db08c08",
  1200 => x"80cf389c",
  1201 => x"160851a7",
  1202 => x"ae2db08c",
  1203 => x"08841b0c",
  1204 => x"9a1680e0",
  1205 => x"2d51a7de",
  1206 => x"2db08c08",
  1207 => x"b08c0888",
  1208 => x"1c0cb08c",
  1209 => x"085555b4",
  1210 => x"fc08802e",
  1211 => x"98389416",
  1212 => x"80e02d51",
  1213 => x"a7de2db0",
  1214 => x"8c08902b",
  1215 => x"83fff00a",
  1216 => x"06701651",
  1217 => x"5473881b",
  1218 => x"0c787a0c",
  1219 => x"7b54a6d2",
  1220 => x"04811858",
  1221 => x"b5800878",
  1222 => x"26fed438",
  1223 => x"b4fc0880",
  1224 => x"2eae387a",
  1225 => x"51a3e42d",
  1226 => x"b08c08b0",
  1227 => x"8c0880ff",
  1228 => x"fffff806",
  1229 => x"555b7380",
  1230 => x"fffffff8",
  1231 => x"2e9238b0",
  1232 => x"8c08fe05",
  1233 => x"b4f40829",
  1234 => x"b5880805",
  1235 => x"57a4e504",
  1236 => x"805473b0",
  1237 => x"8c0c02b4",
  1238 => x"050d0402",
  1239 => x"f4050d74",
  1240 => x"70088105",
  1241 => x"710c7008",
  1242 => x"b4f80806",
  1243 => x"5353718e",
  1244 => x"38881308",
  1245 => x"51a3e42d",
  1246 => x"b08c0888",
  1247 => x"140c810b",
  1248 => x"b08c0c02",
  1249 => x"8c050d04",
  1250 => x"02f0050d",
  1251 => x"75881108",
  1252 => x"fe05b4f4",
  1253 => x"0829b588",
  1254 => x"08117208",
  1255 => x"b4f80806",
  1256 => x"05795553",
  1257 => x"54549bb2",
  1258 => x"2d029005",
  1259 => x"0d0402f4",
  1260 => x"050d7470",
  1261 => x"882a83fe",
  1262 => x"80067072",
  1263 => x"982a0772",
  1264 => x"882b87fc",
  1265 => x"80800673",
  1266 => x"982b81f0",
  1267 => x"0a067173",
  1268 => x"0707b08c",
  1269 => x"0c565153",
  1270 => x"51028c05",
  1271 => x"0d0402f8",
  1272 => x"050d028e",
  1273 => x"0580f52d",
  1274 => x"74882b07",
  1275 => x"7083ffff",
  1276 => x"06b08c0c",
  1277 => x"51028805",
  1278 => x"0d0471b5",
  1279 => x"ac0c0400",
  1280 => x"00ffffff",
  1281 => x"ff00ffff",
  1282 => x"ffff00ff",
  1283 => x"ffffff00",
  1284 => x"20203d20",
  1285 => x"204d5358",
  1286 => x"2d582020",
  1287 => x"203d2020",
  1288 => x"20000000",
  1289 => x"2020204e",
  1290 => x"6575726f",
  1291 => x"52756c65",
  1292 => x"7a202000",
  1293 => x"52657365",
  1294 => x"74000000",
  1295 => x"45786974",
  1296 => x"00000000",
  1297 => x"4b65796d",
  1298 => x"61702045",
  1299 => x"53000000",
  1300 => x"4b65796d",
  1301 => x"61702045",
  1302 => x"4e000000",
  1303 => x"4b65796d",
  1304 => x"61702042",
  1305 => x"52000000",
  1306 => x"4b65796d",
  1307 => x"61702046",
  1308 => x"52000000",
  1309 => x"4f504c33",
  1310 => x"20536f75",
  1311 => x"6e642059",
  1312 => x"65730000",
  1313 => x"4f504c33",
  1314 => x"20536f75",
  1315 => x"6e64204e",
  1316 => x"6f000000",
  1317 => x"52616d20",
  1318 => x"32303438",
  1319 => x"4b420000",
  1320 => x"52616d20",
  1321 => x"34303936",
  1322 => x"4b420000",
  1323 => x"536c6f74",
  1324 => x"20313a20",
  1325 => x"4d656761",
  1326 => x"5343432b",
  1327 => x"20324d42",
  1328 => x"00000000",
  1329 => x"536c6f74",
  1330 => x"20313a20",
  1331 => x"456d7074",
  1332 => x"79536c6f",
  1333 => x"7420313a",
  1334 => x"204d6567",
  1335 => x"6172616d",
  1336 => x"20324d42",
  1337 => x"00000000",
  1338 => x"536c6f74",
  1339 => x"20313a20",
  1340 => x"4d656761",
  1341 => x"72616d20",
  1342 => x"314d4200",
  1343 => x"536c6f74",
  1344 => x"20313a20",
  1345 => x"4d656761",
  1346 => x"5343432b",
  1347 => x"20314d42",
  1348 => x"00000000",
  1349 => x"536c6f74",
  1350 => x"20313a20",
  1351 => x"456d7074",
  1352 => x"79000000",
  1353 => x"536c6f74",
  1354 => x"20303a20",
  1355 => x"45787061",
  1356 => x"6e646564",
  1357 => x"00000000",
  1358 => x"536c6f74",
  1359 => x"20303a20",
  1360 => x"5072696d",
  1361 => x"61727900",
  1362 => x"43505520",
  1363 => x"436c6f63",
  1364 => x"6b204e6f",
  1365 => x"726d616c",
  1366 => x"00000000",
  1367 => x"43505520",
  1368 => x"436c6f63",
  1369 => x"6b205475",
  1370 => x"72626f00",
  1371 => x"426c656e",
  1372 => x"64206f66",
  1373 => x"66000000",
  1374 => x"426c656e",
  1375 => x"64206f6e",
  1376 => x"00000000",
  1377 => x"5363616e",
  1378 => x"6c696e65",
  1379 => x"73204e6f",
  1380 => x"6e650000",
  1381 => x"5363616e",
  1382 => x"6c696e65",
  1383 => x"73204352",
  1384 => x"54203235",
  1385 => x"25000000",
  1386 => x"5363616e",
  1387 => x"6c696e65",
  1388 => x"73204352",
  1389 => x"54203530",
  1390 => x"25000000",
  1391 => x"5363616e",
  1392 => x"6c696e65",
  1393 => x"73204352",
  1394 => x"54203735",
  1395 => x"25000000",
  1396 => x"43617267",
  1397 => x"61204661",
  1398 => x"6c6c6964",
  1399 => x"61000000",
  1400 => x"4f4b0000",
  1401 => x"16200000",
  1402 => x"14200000",
  1403 => x"15200000",
  1404 => x"53442069",
  1405 => x"6e69742e",
  1406 => x"2e2e0a00",
  1407 => x"53442063",
  1408 => x"61726420",
  1409 => x"72657365",
  1410 => x"74206661",
  1411 => x"696c6564",
  1412 => x"210a0000",
  1413 => x"53444843",
  1414 => x"20657272",
  1415 => x"6f72210a",
  1416 => x"00000000",
  1417 => x"57726974",
  1418 => x"65206661",
  1419 => x"696c6564",
  1420 => x"0a000000",
  1421 => x"52656164",
  1422 => x"20666169",
  1423 => x"6c65640a",
  1424 => x"00000000",
  1425 => x"43617264",
  1426 => x"20696e69",
  1427 => x"74206661",
  1428 => x"696c6564",
  1429 => x"0a000000",
  1430 => x"46415431",
  1431 => x"36202020",
  1432 => x"00000000",
  1433 => x"46415433",
  1434 => x"32202020",
  1435 => x"00000000",
  1436 => x"4e6f2070",
  1437 => x"61727469",
  1438 => x"74696f6e",
  1439 => x"20736967",
  1440 => x"0a000000",
  1441 => x"42616420",
  1442 => x"70617274",
  1443 => x"0a000000",
  1444 => x"00000002",
  1445 => x"00000002",
  1446 => x"00001410",
  1447 => x"00000000",
  1448 => x"00000002",
  1449 => x"00001424",
  1450 => x"00000000",
  1451 => x"00000002",
  1452 => x"00001434",
  1453 => x"0000034d",
  1454 => x"00000003",
  1455 => x"00001788",
  1456 => x"00000004",
  1457 => x"00000003",
  1458 => x"00001780",
  1459 => x"00000002",
  1460 => x"00000003",
  1461 => x"00001778",
  1462 => x"00000002",
  1463 => x"00000003",
  1464 => x"00001770",
  1465 => x"00000002",
  1466 => x"00000003",
  1467 => x"00001768",
  1468 => x"00000002",
  1469 => x"00000003",
  1470 => x"0000175c",
  1471 => x"00000004",
  1472 => x"00000003",
  1473 => x"00001754",
  1474 => x"00000002",
  1475 => x"00000003",
  1476 => x"0000174c",
  1477 => x"00000002",
  1478 => x"00000003",
  1479 => x"0000173c",
  1480 => x"00000004",
  1481 => x"00000002",
  1482 => x"0000143c",
  1483 => x"000006e5",
  1484 => x"00000000",
  1485 => x"00000000",
  1486 => x"00000000",
  1487 => x"00001444",
  1488 => x"00001450",
  1489 => x"0000145c",
  1490 => x"00001468",
  1491 => x"00001474",
  1492 => x"00001484",
  1493 => x"00001494",
  1494 => x"000014a0",
  1495 => x"000014ac",
  1496 => x"000014c4",
  1497 => x"000014e8",
  1498 => x"000014fc",
  1499 => x"00001514",
  1500 => x"00001524",
  1501 => x"00001538",
  1502 => x"00001548",
  1503 => x"0000155c",
  1504 => x"0000156c",
  1505 => x"00001578",
  1506 => x"00001584",
  1507 => x"00001594",
  1508 => x"000015a8",
  1509 => x"000015bc",
  1510 => x"00000004",
  1511 => x"000015d0",
  1512 => x"00001798",
  1513 => x"00000004",
  1514 => x"000015e0",
  1515 => x"00001694",
  1516 => x"00000000",
  1517 => x"00000000",
  1518 => x"00000000",
  1519 => x"00000000",
  1520 => x"00000000",
  1521 => x"00000000",
  1522 => x"00000000",
  1523 => x"00000000",
  1524 => x"00000000",
  1525 => x"00000000",
  1526 => x"00000000",
  1527 => x"00000000",
  1528 => x"00000000",
  1529 => x"00000000",
  1530 => x"00000000",
  1531 => x"00000000",
  1532 => x"00000000",
  1533 => x"00000000",
  1534 => x"00000000",
  1535 => x"00000000",
  1536 => x"00000000",
  1537 => x"00000000",
  1538 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

